LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY VGA_display IS
	PORT (
		clock : IN std_logic;
		hcounter : IN INTEGER RANGE 0 TO 1023;
		vcounter : IN INTEGER RANGE 0 TO 1023;
		pixels : OUT std_logic_vector(7 DOWNTO 0)
	);
END VGA_display;

ARCHITECTURE Behavioral OF VGA_display IS
	SIGNAL x : INTEGER RANGE 0 TO 1023 := 100;
	TYPE matrix_type IS ARRAY (0 TO 14, 0 TO 19) OF std_logic_vector(7 DOWNTO 0);
	SIGNAL matrix : matrix_type := (
0=>(0 => B"00000000", 1 => B"00000000", 2 => B"00000000", 3 => B"00000000", 4 => B"00000000", 5=> B"00000000",6=> B"00000000",7=> B"00000000",8=> B"00000000",9=> B"00000000",10=> B"00000000",11=> B"00000000",12=> B"00000000",13=> B"00000000",14=> B"00000000",15=> B"00000000",16=> B"00000000",17=> B"00000000",18=> B"00000000",19=> B"00000000"),
1=>(0 => B"00000000", 1 => B"00000000", 2 => B"00000000", 3 => B"00000000", 4 => B"00000000", 5=> B"00000000",6=> B"00000000",7=> B"00000000",8=> B"00000000",9=> B"00000000",10=> B"00000000",11=> B"00000000",12=> B"00000000",13=> B"00000000",14=> B"00000000",15=> B"00000000",16=> B"00000000",17=> B"00000000",18=> B"00000000",19=> B"00000000"),
2=>(0 => B"00000000", 1 => B"00000000", 2 => B"00000000", 3 => B"00000000", 4 => B"00000000", 5=> B"10010010",6=> B"00000000",7=> B"00000000",8=> B"00000000",9=> B"00000000",10=> B"00000000",11=> B"00000000",12=> B"00000000",13=> B"00000000",14=> B"10010010",15=> B"00000000",16=> B"00000000",17=> B"00000000",18=> B"00000000",19=> B"00000000"),
3=>(0 => B"00000000", 1 => B"00000000", 2 => B"00000000", 3 => B"00000000", 4 => B"00000000", 5=> B"01001001",6=> B"01100000",7=> B"01100000",8=> B"01100000",9=> B"11111111",10=> B"11111111",11=> B"11111111",12=> B"11011011",13=> B"01100000",14=> B"01001001",15=> B"00000000",16=> B"00000000",17=> B"00000000",18=> B"00000000",19=> B"00000000"),
4=>(0 => B"00000000", 1 => B"00000000", 2 => B"00000000", 3 => B"00000000", 4 => B"00000000", 5=> B"01001001",6=> B"01100000",7=> B"01100000",8=> B"01100000",9=> B"11111111",10=> B"11111111",11=> B"11111111",12=> B"01100000",13=> B"01100000",14=> B"01001001",15=> B"00000000",16=> B"00000000",17=> B"00000000",18=> B"00000000",19=> B"00000000"),
5=>(0 => B"00000000", 1 => B"00000000", 2 => B"00000000", 3 => B"00000000", 4 => B"00000000", 5=> B"00000000",6=> B"00000000",7=> B"00000000",8=> B"01100000",9=> B"11111111",10=> B"11111111",11=> B"01100000",12=> B"00000000",13=> B"00000000",14=> B"00000000",15=> B"00000000",16=> B"00000000",17=> B"00000000",18=> B"00000000",19=> B"00000000"),
6=>(0 => B"00000000", 1 => B"00000000", 2 => B"00000000", 3 => B"00000000", 4 => B"00000000", 5=> B"00000000",6=> B"00000000",7=> B"00000000",8=> B"01100000",9=> B"10010010",10=> B"01100000",11=> B"01100000",12=> B"00000000",13=> B"00000000",14=> B"00000000",15=> B"00000000",16=> B"00000000",17=> B"00000000",18=> B"00000000",19=> B"00000000"),
7=>(0 => B"00000000", 1 => B"00000000", 2 => B"00000000", 3 => B"00000000", 4 => B"00000000", 5=> B"00000000",6=> B"01100000",7=> B"01100000",8=> B"01100000",9=> B"01100000",10=> B"01100000",11=> B"01100000",12=> B"01100000",13=> B"01100000",14=> B"00000000",15=> B"00000000",16=> B"00000000",17=> B"00000000",18=> B"00000000",19=> B"00000000"),
8=>(0 => B"00000000", 1 => B"00000000", 2 => B"00000000", 3 => B"00000000", 4 => B"00000000", 5=> B"00000000",6=> B"01100000",7=> B"01100000",8=> B"11111111",9=> B"11111111",10=> B"11111111",11=> B"11111111",12=> B"01100000",13=> B"01100000",14=> B"00000000",15=> B"00000000",16=> B"00000000",17=> B"00000000",18=> B"00000000",19=> B"00000000"),
9=>(0 => B"00000000", 1 => B"00000000", 2 => B"00000000", 3 => B"00000000", 4 => B"00000000", 5=> B"00000000",6=> B"01100000",7=> B"11111111",8=> B"00000000",9=> B"11011011",10=> B"11011011",11=> B"00000000",12=> B"11111111",13=> B"01100000",14=> B"00000000",15=> B"00000000",16=> B"00000000",17=> B"00000000",18=> B"00000000",19=> B"00000000"),
10=>(0 => B"00000000", 1 => B"00000000", 2 => B"00000000", 3 => B"00000000", 4 => B"00000000", 5=> B"00000000",6=> B"01100000",7=> B"11111111",8=> B"11011011",9=> B"10010010",10=> B"10010010",11=> B"11011011",12=> B"11111111",13=> B"01100000",14=> B"00000000",15=> B"00000000",16=> B"00000000",17=> B"00000000",18=> B"00000000",19=> B"00000000"),
11=>(0 => B"00000000", 1 => B"00000000", 2 => B"00000000", 3 => B"00000000", 4 => B"00000000", 5=> B"00000000",6=> B"00000000",7=> B"00000000",8=> B"00000000",9=> B"00000000",10=> B"00000000",11=> B"00000000",12=> B"00000000",13=> B"00000000",14=> B"00000000",15=> B"00000000",16=> B"00000000",17=> B"00000000",18=> B"00000000",19=> B"00000000"),
12=>(0 => B"00000000", 1 => B"00000000", 2 => B"00000000", 3 => B"00000000", 4 => B"00000000", 5=> B"00000000",6=> B"00000000",7=> B"00000000",8=> B"00000000",9=> B"00000000",10=> B"00000000",11=> B"00000000",12=> B"00000000",13=> B"00000000",14=> B"00000000",15=> B"00000000",16=> B"00000000",17=> B"00000000",18=> B"00000000",19=> B"00000000"),
13=>(0 => B"00000000", 1 => B"00000000", 2 => B"00000000", 3 => B"00000000", 4 => B"00000000", 5=> B"00000000",6=> B"00000000",7=> B"00000000",8=> B"00000000",9=> B"00000000",10=> B"00000000",11=> B"00000000",12=> B"00000000",13=> B"00000000",14=> B"00000000",15=> B"00000000",16=> B"00000000",17=> B"00000000",18=> B"00000000",19=> B"00000000"),
14=>(0 => B"00000000", 1 => B"00000000", 2 => B"00000000", 3 => B"00000000", 4 => B"00000000", 5=> B"00000000",6=> B"00000000",7=> B"00000000",8=> B"00000000",9=> B"00000000",10=> B"00000000",11=> B"00000000",12=> B"00000000",13=> B"00000000",14=> B"00000000",15=> B"00000000",16=> B"00000000",17=> B"00000000",18=> B"00000000",19=> B"00000000")
	);
	SIGNAL row_index : INTEGER RANGE 0 TO 14;
	SIGNAL col_index : INTEGER RANGE 0 TO 19;

	-- Constantes
	CONSTANT ROW_DIVISOR : INTEGER := 32;
	CONSTANT COL_DIVISOR : INTEGER := 32;
BEGIN
	video_output : PROCESS (clock)
	BEGIN
		IF rising_edge (clock) THEN
			row_index <= vcounter / ROW_DIVISOR; -- Dividir por 32 para mapear vcounter al rango 0-11
			col_index <= hcounter / COL_DIVISOR; -- Dividir por 32 para mapear hcounter al rango 0-15
			IF (hcounter >= 1) AND (hcounter < 639) AND (vcounter >= 1) AND (vcounter < 479)
			 THEN
			 pixels <= matrix(row_index, col_index);
			 ELSE
				 pixels <= B"00000000";
			 END IF;

		 END IF;
	 END PROCESS;
 END Behavioral;